module logo_table(
		input wire [9:0] addr,
		output wire data
	);

	reg d;
	always @(*) begin
		case (addr)
			0: d = 1'bX;
			1: d = 1'bX;
			2: d = 1'bX;
			3: d = 1'bX;
			4: d = 1'bX;
			5: d = 1'bX;
			6: d = 1'bX;
			7: d = 1'bX;
			8: d = 1'bX;
			9: d = 1'bX;
			10: d = 1'bX;
			11: d = 1'bX;
			12: d = 1'bX;
			13: d = 1'bX;
			14: d = 1'bX;
			15: d = 1'bX;
			16: d = 1'bX;
			17: d = 1'bX;
			18: d = 1'bX;
			19: d = 1'bX;
			20: d = 1'bX;
			21: d = 1'bX;
			22: d = 1'bX;
			23: d = 1'bX;
			24: d = 1'bX;
			25: d = 1'bX;
			26: d = 1'bX;
			27: d = 1'bX;
			28: d = 1'bX;
			29: d = 1'bX;
			30: d = 1'bX;
			31: d = 1'bX;
			32: d = 1'bX;
			33: d = 1'bX;
			34: d = 1'bX;
			35: d = 1'bX;
			36: d = 1'bX;
			37: d = 1'bX;
			38: d = 1'bX;
			39: d = 1'bX;
			40: d = 1'bX;
			41: d = 1'bX;
			42: d = 1'bX;
			43: d = 1'bX;
			44: d = 1'bX;
			45: d = 1'bX;
			46: d = 1'bX;
			47: d = 1'bX;
			48: d = 1'bX;
			49: d = 1'bX;
			50: d = 1'bX;
			51: d = 1'bX;
			52: d = 1'bX;
			53: d = 1'bX;
			54: d = 1'bX;
			55: d = 1'bX;
			56: d = 1'bX;
			57: d = 1'bX;
			58: d = 1'bX;
			59: d = 1'bX;
			60: d = 1'bX;
			61: d = 1'bX;
			62: d = 1'bX;
			63: d = 1'bX;
			64: d = 1'bX;
			65: d = 1'bX;
			66: d = 1'bX;
			67: d = 1'bX;
			68: d = 1'bX;
			69: d = 1'bX;
			70: d = 1'bX;
			71: d = 1'bX;
			72: d = 1'bX;
			73: d = 1'bX;
			74: d = 1'bX;
			75: d = 1'bX;
			76: d = 1'bX;
			77: d = 1'bX;
			78: d = 1'bX;
			79: d = 1'bX;
			80: d = 1'bX;
			81: d = 1'bX;
			82: d = 1'bX;
			83: d = 1'bX;
			84: d = 1'bX;
			85: d = 1'bX;
			86: d = 1'bX;
			87: d = 1'bX;
			88: d = 1'bX;
			89: d = 1'bX;
			90: d = 1'bX;
			91: d = 1'bX;
			92: d = 1'bX;
			93: d = 1'bX;
			94: d = 1'bX;
			95: d = 1'bX;
			96: d = 1'bX;
			97: d = 1'bX;
			98: d = 1'bX;
			99: d = 1'bX;
			100: d = 1'bX;
			101: d = 1'bX;
			102: d = 1'bX;
			103: d = 1'bX;
			104: d = 1'bX;
			105: d = 1'bX;
			106: d = 1'bX;
			107: d = 1'bX;
			108: d = 1'bX;
			109: d = 1'bX;
			110: d = 1'bX;
			111: d = 1'bX;
			112: d = 1'bX;
			113: d = 1'bX;
			114: d = 1'bX;
			115: d = 1'bX;
			116: d = 1'bX;
			117: d = 1'bX;
			118: d = 1'bX;
			119: d = 1'bX;
			120: d = 1'bX;
			121: d = 1'bX;
			122: d = 1'bX;
			123: d = 1'bX;
			124: d = 1'bX;
			125: d = 1'bX;
			126: d = 1'bX;
			127: d = 1'bX;
			128: d = 1'bX;
			129: d = 1'bX;
			130: d = 1'bX;
			131: d = 1'bX;
			132: d = 1'bX;
			133: d = 1'bX;
			134: d = 1'bX;
			135: d = 1'bX;
			136: d = 1'bX;
			137: d = 1'bX;
			138: d = 1'bX;
			139: d = 1'bX;
			140: d = 1'bX;
			141: d = 1'bX;
			142: d = 1'bX;
			143: d = 1'bX;
			144: d = 1'bX;
			145: d = 1'bX;
			146: d = 1'bX;
			147: d = 1'bX;
			148: d = 1'bX;
			149: d = 1'bX;
			150: d = 1'bX;
			151: d = 1'bX;
			152: d = 1'bX;
			153: d = 1'bX;
			154: d = 1'bX;
			155: d = 1'bX;
			156: d = 1'bX;
			157: d = 1'bX;
			158: d = 1'bX;
			159: d = 1'bX;
			160: d = 1'bX;
			161: d = 1'bX;
			162: d = 1'bX;
			163: d = 1'bX;
			164: d = 1'bX;
			165: d = 1'bX;
			166: d = 1'bX;
			167: d = 1'bX;
			168: d = 1'bX;
			169: d = 1'bX;
			170: d = 1'bX;
			171: d = 1'bX;
			172: d = 1'bX;
			173: d = 1'bX;
			174: d = 1'bX;
			175: d = 1'bX;
			176: d = 1'bX;
			177: d = 1'bX;
			178: d = 1'bX;
			179: d = 1'bX;
			180: d = 1'bX;
			181: d = 1'bX;
			182: d = 1'bX;
			183: d = 1'bX;
			184: d = 1'bX;
			185: d = 1'bX;
			186: d = 1'bX;
			187: d = 1'bX;
			188: d = 1'bX;
			189: d = 1'bX;
			190: d = 1'bX;
			191: d = 1'bX;
			192: d = 0;
			193: d = 0;
			194: d = 0;
			195: d = 0;
			196: d = 0;
			197: d = 0;
			198: d = 0;
			199: d = 0;
			200: d = 0;
			201: d = 0;
			202: d = 0;
			203: d = 0;
			204: d = 0;
			205: d = 0;
			206: d = 0;
			207: d = 0;
			208: d = 0;
			209: d = 0;
			210: d = 0;
			211: d = 0;
			212: d = 0;
			213: d = 0;
			214: d = 0;
			215: d = 0;
			216: d = 0;
			217: d = 0;
			218: d = 0;
			219: d = 0;
			220: d = 0;
			221: d = 0;
			222: d = 0;
			223: d = 0;
			224: d = 0;
			225: d = 0;
			226: d = 1;
			227: d = 1;
			228: d = 1;
			229: d = 1;
			230: d = 1;
			231: d = 0;
			232: d = 0;
			233: d = 0;
			234: d = 0;
			235: d = 0;
			236: d = 0;
			237: d = 0;
			238: d = 0;
			239: d = 0;
			240: d = 0;
			241: d = 0;
			242: d = 0;
			243: d = 0;
			244: d = 0;
			245: d = 0;
			246: d = 0;
			247: d = 0;
			248: d = 0;
			249: d = 0;
			250: d = 0;
			251: d = 0;
			252: d = 0;
			253: d = 0;
			254: d = 0;
			255: d = 0;
			256: d = 0;
			257: d = 0;
			258: d = 1;
			259: d = 1;
			260: d = 1;
			261: d = 0;
			262: d = 1;
			263: d = 1;
			264: d = 0;
			265: d = 0;
			266: d = 0;
			267: d = 0;
			268: d = 0;
			269: d = 0;
			270: d = 0;
			271: d = 0;
			272: d = 0;
			273: d = 0;
			274: d = 0;
			275: d = 0;
			276: d = 0;
			277: d = 0;
			278: d = 0;
			279: d = 0;
			280: d = 0;
			281: d = 0;
			282: d = 0;
			283: d = 0;
			284: d = 0;
			285: d = 0;
			286: d = 0;
			287: d = 0;
			288: d = 0;
			289: d = 0;
			290: d = 0;
			291: d = 1;
			292: d = 1;
			293: d = 1;
			294: d = 1;
			295: d = 1;
			296: d = 0;
			297: d = 0;
			298: d = 0;
			299: d = 0;
			300: d = 0;
			301: d = 0;
			302: d = 0;
			303: d = 0;
			304: d = 0;
			305: d = 0;
			306: d = 0;
			307: d = 0;
			308: d = 0;
			309: d = 0;
			310: d = 0;
			311: d = 0;
			312: d = 0;
			313: d = 0;
			314: d = 0;
			315: d = 0;
			316: d = 0;
			317: d = 0;
			318: d = 0;
			319: d = 0;
			320: d = 0;
			321: d = 0;
			322: d = 0;
			323: d = 0;
			324: d = 0;
			325: d = 0;
			326: d = 0;
			327: d = 0;
			328: d = 0;
			329: d = 0;
			330: d = 0;
			331: d = 1;
			332: d = 1;
			333: d = 1;
			334: d = 1;
			335: d = 1;
			336: d = 0;
			337: d = 0;
			338: d = 0;
			339: d = 0;
			340: d = 0;
			341: d = 0;
			342: d = 0;
			343: d = 0;
			344: d = 0;
			345: d = 0;
			346: d = 0;
			347: d = 0;
			348: d = 0;
			349: d = 0;
			350: d = 0;
			351: d = 0;
			352: d = 0;
			353: d = 0;
			354: d = 1;
			355: d = 1;
			356: d = 1;
			357: d = 1;
			358: d = 1;
			359: d = 1;
			360: d = 0;
			361: d = 0;
			362: d = 0;
			363: d = 0;
			364: d = 0;
			365: d = 0;
			366: d = 0;
			367: d = 0;
			368: d = 0;
			369: d = 0;
			370: d = 0;
			371: d = 0;
			372: d = 0;
			373: d = 0;
			374: d = 0;
			375: d = 0;
			376: d = 0;
			377: d = 0;
			378: d = 0;
			379: d = 0;
			380: d = 0;
			381: d = 0;
			382: d = 0;
			383: d = 0;
			384: d = 0;
			385: d = 0;
			386: d = 1;
			387: d = 1;
			388: d = 1;
			389: d = 0;
			390: d = 1;
			391: d = 0;
			392: d = 0;
			393: d = 0;
			394: d = 1;
			395: d = 1;
			396: d = 1;
			397: d = 1;
			398: d = 1;
			399: d = 1;
			400: d = 0;
			401: d = 0;
			402: d = 0;
			403: d = 0;
			404: d = 0;
			405: d = 0;
			406: d = 0;
			407: d = 0;
			408: d = 0;
			409: d = 0;
			410: d = 0;
			411: d = 0;
			412: d = 0;
			413: d = 0;
			414: d = 0;
			415: d = 0;
			416: d = 0;
			417: d = 0;
			418: d = 0;
			419: d = 1;
			420: d = 1;
			421: d = 1;
			422: d = 0;
			423: d = 1;
			424: d = 0;
			425: d = 0;
			426: d = 1;
			427: d = 1;
			428: d = 1;
			429: d = 0;
			430: d = 1;
			431: d = 0;
			432: d = 0;
			433: d = 0;
			434: d = 0;
			435: d = 0;
			436: d = 0;
			437: d = 0;
			438: d = 0;
			439: d = 0;
			440: d = 0;
			441: d = 0;
			442: d = 0;
			443: d = 0;
			444: d = 0;
			445: d = 0;
			446: d = 0;
			447: d = 0;
			448: d = 0;
			449: d = 0;
			450: d = 0;
			451: d = 0;
			452: d = 0;
			453: d = 0;
			454: d = 0;
			455: d = 0;
			456: d = 0;
			457: d = 0;
			458: d = 0;
			459: d = 1;
			460: d = 1;
			461: d = 1;
			462: d = 0;
			463: d = 1;
			464: d = 0;
			465: d = 0;
			466: d = 0;
			467: d = 0;
			468: d = 0;
			469: d = 0;
			470: d = 0;
			471: d = 0;
			472: d = 0;
			473: d = 0;
			474: d = 0;
			475: d = 0;
			476: d = 0;
			477: d = 0;
			478: d = 0;
			479: d = 0;
			480: d = 0;
			481: d = 0;
			482: d = 0;
			483: d = 1;
			484: d = 1;
			485: d = 1;
			486: d = 1;
			487: d = 1;
			488: d = 0;
			489: d = 0;
			490: d = 0;
			491: d = 0;
			492: d = 0;
			493: d = 0;
			494: d = 0;
			495: d = 0;
			496: d = 0;
			497: d = 0;
			498: d = 0;
			499: d = 1;
			500: d = 1;
			501: d = 1;
			502: d = 1;
			503: d = 1;
			504: d = 0;
			505: d = 0;
			506: d = 0;
			507: d = 0;
			508: d = 0;
			509: d = 0;
			510: d = 0;
			511: d = 0;
			512: d = 0;
			513: d = 0;
			514: d = 0;
			515: d = 0;
			516: d = 0;
			517: d = 0;
			518: d = 0;
			519: d = 0;
			520: d = 0;
			521: d = 0;
			522: d = 1;
			523: d = 1;
			524: d = 1;
			525: d = 1;
			526: d = 1;
			527: d = 0;
			528: d = 0;
			529: d = 0;
			530: d = 0;
			531: d = 0;
			532: d = 0;
			533: d = 0;
			534: d = 0;
			535: d = 0;
			536: d = 0;
			537: d = 0;
			538: d = 0;
			539: d = 0;
			540: d = 0;
			541: d = 0;
			542: d = 0;
			543: d = 0;
			544: d = 0;
			545: d = 0;
			546: d = 1;
			547: d = 1;
			548: d = 1;
			549: d = 1;
			550: d = 1;
			551: d = 0;
			552: d = 0;
			553: d = 0;
			554: d = 1;
			555: d = 1;
			556: d = 1;
			557: d = 0;
			558: d = 1;
			559: d = 1;
			560: d = 0;
			561: d = 0;
			562: d = 1;
			563: d = 1;
			564: d = 1;
			565: d = 1;
			566: d = 1;
			567: d = 0;
			568: d = 0;
			569: d = 0;
			570: d = 1;
			571: d = 1;
			572: d = 1;
			573: d = 1;
			574: d = 1;
			575: d = 0;
			576: d = 0;
			577: d = 0;
			578: d = 1;
			579: d = 1;
			580: d = 1;
			581: d = 0;
			582: d = 1;
			583: d = 1;
			584: d = 0;
			585: d = 0;
			586: d = 0;
			587: d = 1;
			588: d = 1;
			589: d = 1;
			590: d = 1;
			591: d = 1;
			592: d = 0;
			593: d = 0;
			594: d = 1;
			595: d = 1;
			596: d = 1;
			597: d = 0;
			598: d = 1;
			599: d = 1;
			600: d = 0;
			601: d = 0;
			602: d = 1;
			603: d = 1;
			604: d = 1;
			605: d = 0;
			606: d = 1;
			607: d = 1;
			608: d = 0;
			609: d = 0;
			610: d = 0;
			611: d = 1;
			612: d = 1;
			613: d = 1;
			614: d = 1;
			615: d = 1;
			616: d = 0;
			617: d = 0;
			618: d = 0;
			619: d = 0;
			620: d = 0;
			621: d = 0;
			622: d = 0;
			623: d = 0;
			624: d = 0;
			625: d = 0;
			626: d = 0;
			627: d = 1;
			628: d = 1;
			629: d = 1;
			630: d = 1;
			631: d = 1;
			632: d = 0;
			633: d = 0;
			634: d = 0;
			635: d = 1;
			636: d = 1;
			637: d = 1;
			638: d = 1;
			639: d = 1;
			640: d = 0;
			641: d = 0;
			642: d = 0;
			643: d = 0;
			644: d = 0;
			645: d = 0;
			646: d = 0;
			647: d = 0;
			648: d = 0;
			649: d = 0;
			650: d = 1;
			651: d = 1;
			652: d = 1;
			653: d = 1;
			654: d = 1;
			655: d = 1;
			656: d = 0;
			657: d = 0;
			658: d = 0;
			659: d = 0;
			660: d = 0;
			661: d = 0;
			662: d = 0;
			663: d = 0;
			664: d = 0;
			665: d = 0;
			666: d = 0;
			667: d = 0;
			668: d = 0;
			669: d = 0;
			670: d = 0;
			671: d = 0;
			672: d = 0;
			673: d = 0;
			674: d = 1;
			675: d = 1;
			676: d = 1;
			677: d = 1;
			678: d = 1;
			679: d = 1;
			680: d = 0;
			681: d = 0;
			682: d = 0;
			683: d = 1;
			684: d = 1;
			685: d = 1;
			686: d = 1;
			687: d = 0;
			688: d = 0;
			689: d = 0;
			690: d = 1;
			691: d = 1;
			692: d = 1;
			693: d = 1;
			694: d = 1;
			695: d = 1;
			696: d = 0;
			697: d = 0;
			698: d = 1;
			699: d = 1;
			700: d = 1;
			701: d = 1;
			702: d = 1;
			703: d = 1;
			704: d = 0;
			705: d = 0;
			706: d = 0;
			707: d = 1;
			708: d = 1;
			709: d = 1;
			710: d = 1;
			711: d = 0;
			712: d = 0;
			713: d = 0;
			714: d = 0;
			715: d = 1;
			716: d = 1;
			717: d = 1;
			718: d = 1;
			719: d = 1;
			720: d = 0;
			721: d = 0;
			722: d = 0;
			723: d = 1;
			724: d = 1;
			725: d = 1;
			726: d = 1;
			727: d = 0;
			728: d = 0;
			729: d = 0;
			730: d = 0;
			731: d = 1;
			732: d = 1;
			733: d = 1;
			734: d = 1;
			735: d = 0;
			736: d = 0;
			737: d = 0;
			738: d = 0;
			739: d = 1;
			740: d = 1;
			741: d = 1;
			742: d = 1;
			743: d = 1;
			744: d = 0;
			745: d = 0;
			746: d = 0;
			747: d = 0;
			748: d = 0;
			749: d = 0;
			750: d = 0;
			751: d = 0;
			752: d = 0;
			753: d = 0;
			754: d = 0;
			755: d = 1;
			756: d = 1;
			757: d = 1;
			758: d = 1;
			759: d = 1;
			760: d = 0;
			761: d = 0;
			762: d = 0;
			763: d = 1;
			764: d = 1;
			765: d = 1;
			766: d = 1;
			767: d = 1;
			768: d = 0;
			769: d = 0;
			770: d = 0;
			771: d = 0;
			772: d = 0;
			773: d = 0;
			774: d = 0;
			775: d = 0;
			776: d = 0;
			777: d = 0;
			778: d = 0;
			779: d = 0;
			780: d = 0;
			781: d = 0;
			782: d = 0;
			783: d = 0;
			784: d = 0;
			785: d = 0;
			786: d = 0;
			787: d = 0;
			788: d = 0;
			789: d = 0;
			790: d = 0;
			791: d = 0;
			792: d = 0;
			793: d = 0;
			794: d = 0;
			795: d = 0;
			796: d = 0;
			797: d = 0;
			798: d = 0;
			799: d = 0;
			800: d = 0;
			801: d = 0;
			802: d = 0;
			803: d = 0;
			804: d = 0;
			805: d = 0;
			806: d = 0;
			807: d = 0;
			808: d = 0;
			809: d = 0;
			810: d = 0;
			811: d = 0;
			812: d = 0;
			813: d = 0;
			814: d = 0;
			815: d = 0;
			816: d = 0;
			817: d = 0;
			818: d = 0;
			819: d = 0;
			820: d = 0;
			821: d = 0;
			822: d = 0;
			823: d = 0;
			824: d = 0;
			825: d = 0;
			826: d = 0;
			827: d = 0;
			828: d = 0;
			829: d = 0;
			830: d = 0;
			831: d = 0;
			832: d = 1'bX;
			833: d = 1'bX;
			834: d = 1'bX;
			835: d = 1'bX;
			836: d = 1'bX;
			837: d = 1'bX;
			838: d = 1'bX;
			839: d = 1'bX;
			840: d = 1'bX;
			841: d = 1'bX;
			842: d = 1'bX;
			843: d = 1'bX;
			844: d = 1'bX;
			845: d = 1'bX;
			846: d = 1'bX;
			847: d = 1'bX;
			848: d = 1'bX;
			849: d = 1'bX;
			850: d = 1'bX;
			851: d = 1'bX;
			852: d = 1'bX;
			853: d = 1'bX;
			854: d = 1'bX;
			855: d = 1'bX;
			856: d = 1'bX;
			857: d = 1'bX;
			858: d = 1'bX;
			859: d = 1'bX;
			860: d = 1'bX;
			861: d = 1'bX;
			862: d = 1'bX;
			863: d = 1'bX;
			864: d = 1'bX;
			865: d = 1'bX;
			866: d = 1'bX;
			867: d = 1'bX;
			868: d = 1'bX;
			869: d = 1'bX;
			870: d = 1'bX;
			871: d = 1'bX;
			872: d = 1'bX;
			873: d = 1'bX;
			874: d = 1'bX;
			875: d = 1'bX;
			876: d = 1'bX;
			877: d = 1'bX;
			878: d = 1'bX;
			879: d = 1'bX;
			880: d = 1'bX;
			881: d = 1'bX;
			882: d = 1'bX;
			883: d = 1'bX;
			884: d = 1'bX;
			885: d = 1'bX;
			886: d = 1'bX;
			887: d = 1'bX;
			888: d = 1'bX;
			889: d = 1'bX;
			890: d = 1'bX;
			891: d = 1'bX;
			892: d = 1'bX;
			893: d = 1'bX;
			894: d = 1'bX;
			895: d = 1'bX;
			896: d = 1'bX;
			897: d = 1'bX;
			898: d = 1'bX;
			899: d = 1'bX;
			900: d = 1'bX;
			901: d = 1'bX;
			902: d = 1'bX;
			903: d = 1'bX;
			904: d = 1'bX;
			905: d = 1'bX;
			906: d = 1'bX;
			907: d = 1'bX;
			908: d = 1'bX;
			909: d = 1'bX;
			910: d = 1'bX;
			911: d = 1'bX;
			912: d = 1'bX;
			913: d = 1'bX;
			914: d = 1'bX;
			915: d = 1'bX;
			916: d = 1'bX;
			917: d = 1'bX;
			918: d = 1'bX;
			919: d = 1'bX;
			920: d = 1'bX;
			921: d = 1'bX;
			922: d = 1'bX;
			923: d = 1'bX;
			924: d = 1'bX;
			925: d = 1'bX;
			926: d = 1'bX;
			927: d = 1'bX;
			928: d = 1'bX;
			929: d = 1'bX;
			930: d = 1'bX;
			931: d = 1'bX;
			932: d = 1'bX;
			933: d = 1'bX;
			934: d = 1'bX;
			935: d = 1'bX;
			936: d = 1'bX;
			937: d = 1'bX;
			938: d = 1'bX;
			939: d = 1'bX;
			940: d = 1'bX;
			941: d = 1'bX;
			942: d = 1'bX;
			943: d = 1'bX;
			944: d = 1'bX;
			945: d = 1'bX;
			946: d = 1'bX;
			947: d = 1'bX;
			948: d = 1'bX;
			949: d = 1'bX;
			950: d = 1'bX;
			951: d = 1'bX;
			952: d = 1'bX;
			953: d = 1'bX;
			954: d = 1'bX;
			955: d = 1'bX;
			956: d = 1'bX;
			957: d = 1'bX;
			958: d = 1'bX;
			959: d = 1'bX;
			960: d = 1'bX;
			961: d = 1'bX;
			962: d = 1'bX;
			963: d = 1'bX;
			964: d = 1'bX;
			965: d = 1'bX;
			966: d = 1'bX;
			967: d = 1'bX;
			968: d = 1'bX;
			969: d = 1'bX;
			970: d = 1'bX;
			971: d = 1'bX;
			972: d = 1'bX;
			973: d = 1'bX;
			974: d = 1'bX;
			975: d = 1'bX;
			976: d = 1'bX;
			977: d = 1'bX;
			978: d = 1'bX;
			979: d = 1'bX;
			980: d = 1'bX;
			981: d = 1'bX;
			982: d = 1'bX;
			983: d = 1'bX;
			984: d = 1'bX;
			985: d = 1'bX;
			986: d = 1'bX;
			987: d = 1'bX;
			988: d = 1'bX;
			989: d = 1'bX;
			990: d = 1'bX;
			991: d = 1'bX;
			992: d = 1'bX;
			993: d = 1'bX;
			994: d = 1'bX;
			995: d = 1'bX;
			996: d = 1'bX;
			997: d = 1'bX;
			998: d = 1'bX;
			999: d = 1'bX;
			1000: d = 1'bX;
			1001: d = 1'bX;
			1002: d = 1'bX;
			1003: d = 1'bX;
			1004: d = 1'bX;
			1005: d = 1'bX;
			1006: d = 1'bX;
			1007: d = 1'bX;
			1008: d = 1'bX;
			1009: d = 1'bX;
			1010: d = 1'bX;
			1011: d = 1'bX;
			1012: d = 1'bX;
			1013: d = 1'bX;
			1014: d = 1'bX;
			1015: d = 1'bX;
			1016: d = 1'bX;
			1017: d = 1'bX;
			1018: d = 1'bX;
			1019: d = 1'bX;
			1020: d = 1'bX;
			1021: d = 1'bX;
			1022: d = 1'bX;
			1023: d = 1'bX;
			default: d = 'X;
		endcase
	end

	assign data = d;
endmodule : logo_table
