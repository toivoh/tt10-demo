/*
 * Copyright (c) 2025 Toivo Henningsson
 * SPDX-License-Identifier: Apache-2.0
 */

`define DEMO_TIME_BITS 13

`ifndef FPGA
`define DEMO_TIME_START 512
//`define DEMO_TIME_START (5*1024 + 4*8)
`else
`define DEMO_TIME_START 512
//`define DEMO_TIME_START (2*1024 - 256)
//`define DEMO_TIME_START (3*1024 - 256)
//`define DEMO_TIME_START (4*1024 - 256)
//`define DEMO_TIME_START (6*1024 - 256)
`endif

`define PATTERN_BITS 2

`define AFL_SECTION_BITS 1
`define AFL_SECTION_PILLAR 1'd0
`define AFL_SECTION_SPIRAL 1'd1
/*
`define AFL_SECTION_BITS 2
`define AFL_SECTION_PILLAR 2'd0
`define AFL_SECTION_SPIRAL 2'd1
`define AFL_SECTION_RP     2'd2
*/

`define WAVE_MODE_BITS 2
`define WAVE_MODE_PRENOISE 2'd0
`define WAVE_MODE_BASS     2'd1
`define WAVE_MODE_DRUMS    2'd2
`define WAVE_MODE_ARP      2'd3


`define DEMO_CONTROL_BIT_MELODY 0
`define DEMO_CONTROL_BIT_BDRUM 1
`define DEMO_CONTROL_BIT_NDRUM 2
`define DEMO_CONTROL_BIT_BASS 3
`define DEMO_CONTROL_BIT_NOISE 4
`define DEMO_CONTROL_BIT_RAISE 5
`define DEMO_CONTROL_BIT_PRENOISE 6
`define DEMO_CONTROL_BIT_SQUARE 7
`define DEMO_CONTROL_BIT_EFFECT 8
`define DEMO_CONTROL_BIT_DETUNE_DOUBLE 9
`define DEMO_CONTROL_BIT_LOGO_ON 10
`define DEMO_CONTROL_BIT_LOGO_LINES0 11
`define DEMO_CONTROL_BIT_LOGO_LINES1 12
`define DEMO_CONTROL_BIT_REV_LOGO_LINES 13
`define DEMO_CONTROL_BIT_WAVE_ON 14

`define DEMO_CONTROL_BIT_PATTERN 15
`define DEMO_CONTROL_BIT_AFL (`DEMO_CONTROL_BIT_PATTERN + `PATTERN_BITS)
`define DEMO_CONTROL_BIT_WAVE_MODE (`DEMO_CONTROL_BIT_PATTERN + `PATTERN_BITS + `AFL_SECTION_BITS)
`define DEMO_CONTROL_BITS (`DEMO_CONTROL_BIT_PATTERN + `PATTERN_BITS + `AFL_SECTION_BITS + `WAVE_MODE_BITS)


//`define DEBUG_ON
//`define SMALL


`ifdef SMALL
//`define USE_FIELD

//`define OSC_BITS 21
//`define POS_BITS 7
//`define POS_BITS_GT1_PATTERN

`define OSC_BITS 22
`define POS_BITS 9
`define POS_BITS_GT1_PATTERN
`else
`define USE_FIELD
`define USE_AFL
`define USE_LOGO
`define OSC_BITS 23
`define POS_BITS 9
`define POS_BITS_GT1_PATTERN
`endif


`define USE_AFL_MC
`define USE_RAISE
`define USE_SEMITONE_CODING

`ifdef USE_RAISE
`define USE_SEMITONE_CODING
`endif
